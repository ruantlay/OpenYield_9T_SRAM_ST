* 9T SRAM RSNM - Xyce Compatibility Fix
.INCLUDE "tmp_mc.spice"

* --- 电源定义 ---
VVDD VDD 0 0.5
VVSS VSS 0 0
VWL  WL  0 0.5
VBL  BL  0 0.5
VWWLA WWLA 0 0
VWWLB WWLB_NET 0 0.5
VSCAN VIN_COMMON 0 0

* --- 9T 电路结构 ---
* 左侧支路
MPUL1  V1  VIN_COMMON VDD VDD PMOS_VTG W=120n L=60n
MPUL2  VQ  WWLA       V1  VDD PMOS_VTG W=120n L=60n
MNPDL1 VQ  VDD        V2  VSS NMOS_VTG W=100n L=60n 
MNPDL2 V2  VIN_COMMON VSS VSS NMOS_VTG W=100n L=60n
MPG    VQ  WL         BL  VSS NMOS_VTG W=60n  L=50n

* 右侧 ST 结构 (根据论文, MNF 决定迟滞特性)
MPUR  VQB VIN_COMMON VDD VDD PMOS_VTG W=120n L=150n
MPDR1 VQB VIN_COMMON VX  VSS NMOS_VTG W=80n  L=60n
MPDR2 VX  VIN_COMMON VSS VSS NMOS_VTG W=80n  L=60n
MNF   VX  VQB WWLB_NET VSS NMOS_VTG W=40n  L=100n

* --- 修正后的 DC 扫描语句 ---
* Xyce 双重扫描语法格式：.DC 变量1 起始 终止 步长 变量2 起始 终止 步长
.DC VSCAN 0 0.5 0.005 VWWLB 0.3 0.5 0.1

* 导出数据
.PRINT DC FORMAT=CSV FILE=RSNM_DATA.csv V(VIN_COMMON) V(VQ) V(VQB) V(WWLB_NET)
.END