.model  NMOS_VTL  nmos
+       level = 54                                tnom = 27                              epsrox = 3.9                               eta0 = 0.006                     
+     nfactor = 2.1                               wint = 5.000e-09                         cgso = 1.100e-10                         cgdo = 1.100e-10                 
+          xl = -2.000e-08                        toxe = 1.140e-09                         toxp = 1.000e-09                         toxm = 1.140e-09                 
+      toxref = 1.140e-09                         dtox = 1.400e-10                         lint = 3.750e-09                         vth0 = {AGAUSS(0.322, 0.01610, 1)}
+          k1 = 0.4                                 u0 = {AGAUSS(0.045, 0.00225, 1)}        vsat = 148000                            rdsw = 155                       
+        ndep = 3.400e+18                           xj = 1.980e-08                      version = 4.8                            binunit = 1                         
+    paramchk = 1                               mobmod = 0                               capmod = 2                               igcmod = 1                         
+      igbmod = 1                               geomod = 1                               diomod = 1                               rdsmod = 0                         
+    rbodymod = 1                             rgatemod = 1                               permod = 1                             acnqsmod = 0                         
+    trnqsmod = 0                                   ll = 0                                   wl = 0                                  lln = 1                         
+         wln = 1                                   lw = 0                                   ww = 0                                  lwn = 1                         
+         wwn = 1                                  lwl = 0                                  wwl = 0                                xpart = 0                         
+          k2 = 0                                   k3 = 0                                  k3b = 0                                   w0 = 2.500e-06                 
+        dvt0 = 1                                 dvt1 = 2                                 dvt2 = 0                                dvt0w = 0                         
+       dvt1w = 0                                dvt2w = 0                                 dsub = 0.1                               minv = 0.05                      
+       voffl = 0                                dvtp0 = 1.000e-10                        dvtp1 = 0.1                               lpe0 = 0                         
+        lpeb = 0                                ngate = 3.000e+20                          nsd = 2.000e+20                         phin = 0                         
+        cdsc = 0                                cdscb = 0                                cdscd = 0                                  cit = 0                         
+        voff = {AGAUSS(-0.13, 0.00650, 1)}        etab = 0                                  vfb = -0.55                               ua = 6.000e-10                 
+          ub = 1.200e-18                           uc = 0                                   a0 = 1                                  ags = 0                         
+          a1 = 0                                   a2 = 1                                   b0 = 0                                   b1 = 0                         
+        keta = 0.04                               dwg = 0                                  dwb = 0                                 pclm = 0.02                      
+     pdiblc1 = 0.001                          pdiblc2 = 0.001                          pdiblcb = -0.005                           drout = 0.5                       
+        pvag = 1.000e-20                        delta = 0.01                            pscbe1 = 8.140e+08                       pscbe2 = 1.000e-07                 
+      fprout = 0.2                              pdits = 0.08                            pditsd = 0.23                            pditsl = 2300000                   
+         rsh = 5                                  rsw = 80                                 rdw = 80                             rdswmin = 0                         
+      rdwmin = 0                               rswmin = 0                                 prwg = 0                                 prwb = 0                         
+          wr = 1                               alpha0 = 0.074                           alpha1 = 0.005                            beta0 = 30                        
+       agidl = 2.000e-04                        bgidl = 2.100e+09                        cgidl = 2.000e-04                        egidl = 0.8                       
+     aigbacc = 0.012                          bigbacc = 0.0028                         cigbacc = 0.002                          nigbacc = 1                         
+     aigbinv = 0.014                          bigbinv = 0.004                          cigbinv = 0.004                          eigbinv = 1.1                       
+     nigbinv = 3                                 aigc = 0.02                              bigc = 0.0027                            cigc = 0.002                     
+       aigsd = 0.02                             bigsd = 0.0027                           cigsd = 0.002                             nigc = 1                         
+     poxedge = 1                                pigcd = 1                                 ntox = 1                               xrcrg1 = 12                        
+      xrcrg2 = 5                                 cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                 
+     ckappas = 0.03                           ckappad = 0.03                              acde = 1                                 moin = 15                        
+        noff = 0.9                             voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                         
+         kt2 = 0.022                              ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                 
+         uc1 = -5.600e-11                         prt = 0                                   at = 33000                          fnoimod = 1                         
+     tnoimod = 0                                  jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                 
+         njs = 1                             ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                        
+       xjbvs = 1                                  jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                 
+         njd = 1                             ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                        
+       xjbvd = 1                                  pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                       
+       pbsws = 1                                cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                         
+      cjswgs = 3.000e-10                       mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                 
+         mjd = 0.5                              pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                      
+      pbswgd = 1                               cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                     
+         tcj = 0.001                            tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                     
+      tcjswg = 0.001                             xtis = 3                                 xtid = 3                                 dmcg = 0                         
+        dmci = 0                                 dmdg = 0                                dmcgt = 0                                  dwj = 0                         
+         xgw = 0                                  xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                 
+        rbpb = 5                                 rbpd = 15                                rbps = 15                                rbdb = 15                        
+        rbsb = 15                               ngcon = 1                         

.model  PMOS_VTL  pmos
+       level = 54                                vth0 = {AGAUSS(-0.3021, 0.01511, 1)}      toxref = 1.300e-09                         vsat = 69000                     
+        toxe = 1.260e-09                         toxp = 1.000e-09                         toxm = 1.260e-09                         dtox = 2.600e-10                 
+      epsrox = 3.9                               wint = 5.000e-09                         lint = 3.750e-09                      version = 4.8                       
+     binunit = 1                             paramchk = 1                               mobmod = 0                               capmod = 2                         
+      igcmod = 1                               igbmod = 1                               geomod = 1                               diomod = 1                         
+      rdsmod = 0                             rbodymod = 1                             rgatemod = 1                               permod = 1                         
+    acnqsmod = 0                             trnqsmod = 0                                 tnom = 27                                  ll = 0                         
+          wl = 0                                  lln = 1                                  wln = 1                                   lw = 0                         
+          ww = 0                                  lwn = 1                                  wwn = 1                                  lwl = 0                         
+         wwl = 0                                xpart = 0                                   xl = -2.000e-08                          k1 = 0.4                       
+          k2 = -0.01                               k3 = 0                                  k3b = 0                                   w0 = 2.500e-06                 
+        dvt0 = 1                                 dvt1 = 2                                 dvt2 = -0.032                           dvt0w = 0                         
+       dvt1w = 0                                dvt2w = 0                                 dsub = 0.1                               minv = 0.05                      
+       voffl = 0                                dvtp0 = 1.000e-11                        dvtp1 = 0.05                              lpe0 = 0                         
+        lpeb = 0                                   xj = 1.980e-08                        ngate = 2.000e+20                         ndep = 2.440e+18                 
+         nsd = 2.000e+20                         phin = 0                                 cdsc = 0                                cdscb = 0                         
+       cdscd = 0                                  cit = 0                                 voff = {AGAUSS(-0.126, 0.00630, 1)}     nfactor = 2.22                      
+        eta0 = 0.0055                            etab = 0                                  vfb = 0.55                                u0 = {AGAUSS(0.02, 0.00100, 1)}
+          ua = 2.000e-09                           ub = 5.000e-19                           uc = 0                                   a0 = 1                         
+         ags = 1.000e-20                           a1 = 0                                   a2 = 1                                   b0 = 0                         
+          b1 = 0                                 keta = -0.047                             dwg = 0                                  dwb = 0                         
+        pclm = 0.12                           pdiblc1 = 0.001                          pdiblc2 = 0.001                          pdiblcb = 3.400e-08                 
+       drout = 0.56                              pvag = 1.000e-20                        delta = 0.01                            pscbe1 = 8.140e+08                 
+      pscbe2 = 9.580e-07                       fprout = 0.2                              pdits = 0.08                            pditsd = 0.23                      
+      pditsl = 2300000                            rsh = 5                                 rdsw = 155                                rsw = 75                        
+         rdw = 75                             rdswmin = 0                               rdwmin = 0                               rswmin = 0                         
+        prwg = 0                                 prwb = 0                                   wr = 1                               alpha0 = 0.074                     
+      alpha1 = 0.005                            beta0 = 30                               agidl = 2.000e-04                        bgidl = 2.100e+09                 
+       cgidl = 2.000e-04                        egidl = 0.8                            aigbacc = 0.012                          bigbacc = 0.0028                    
+     cigbacc = 0.002                          nigbacc = 1                              aigbinv = 0.014                          bigbinv = 0.004                     
+     cigbinv = 0.004                          eigbinv = 1.1                            nigbinv = 3                                 aigc = 0.010687                  
+        bigc = 0.0012607                         cigc = 8.000e-04                        aigsd = 0.010687                         bigsd = 0.0012607                 
+       cigsd = 8.000e-04                         nigc = 1                              poxedge = 1                                pigcd = 1                         
+        ntox = 1                               xrcrg1 = 12                              xrcrg2 = 5                                 cgso = 1.100e-10                 
+        cgdo = 1.100e-10                         cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                 
+     ckappas = 0.03                           ckappad = 0.03                              acde = 1                                 moin = 15                        
+        noff = 0.9                             voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                         
+         kt2 = 0.022                              ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                 
+         uc1 = -5.600e-11                         prt = 0                                   at = 33000                          fnoimod = 1                         
+     tnoimod = 0                                  jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                 
+         njs = 1                             ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                        
+       xjbvs = 1                                  jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                 
+         njd = 1                             ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                        
+       xjbvd = 1                                  pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                       
+       pbsws = 1                                cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                         
+      cjswgs = 3.000e-10                       mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                 
+         mjd = 0.5                              pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                      
+      pbswgd = 1                               cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                     
+         tcj = 0.001                            tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                     
+      tcjswg = 0.001                             xtis = 3                                 xtid = 3                                 dmcg = 0                         
+        dmci = 0                                 dmdg = 0                                dmcgt = 0                                  dwj = 0                         
+         xgw = 0                                  xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                 
+        rbpb = 5                                 rbpd = 15                                rbps = 15                                rbdb = 15                        
+        rbsb = 15                               ngcon = 1                         

.model  NMOS_VTG  nmos
+       level = 54                                tnom = 27                              epsrox = 3.9                               eta0 = 0.006                     
+     nfactor = 2.1                               wint = 5.000e-09                         cgso = 1.100e-10                         cgdo = 1.100e-10                 
+          xl = -2.000e-08                        toxe = 1.140e-09                         toxp = 1.000e-09                         toxm = 1.140e-09                 
+      toxref = 1.140e-09                         dtox = 1.400e-10                         lint = 3.750e-09                         vth0 = {AGAUSS(0.4106, 0.02053, 1)}
+          k1 = 0.4                                 u0 = {AGAUSS(0.045, 0.00225, 1)}        vsat = 123000                            rdsw = 155                       
+        ndep = 3.400e+18                           xj = 1.980e-08                      version = 4.8                            binunit = 1                         
+    paramchk = 1                               mobmod = 0                               capmod = 2                               igcmod = 1                         
+      igbmod = 1                               geomod = 1                               diomod = 1                               rdsmod = 0                         
+    rbodymod = 1                             rgatemod = 1                               permod = 1                             acnqsmod = 0                         
+    trnqsmod = 0                                   ll = 0                                   wl = 0                                  lln = 1                         
+         wln = 1                                   lw = 0                                   ww = 0                                  lwn = 1                         
+         wwn = 1                                  lwl = 0                                  wwl = 0                                xpart = 0                         
+          k2 = 0                                   k3 = 0                                  k3b = 0                                   w0 = 2.500e-06                 
+        dvt0 = 1                                 dvt1 = 2                                 dvt2 = 0                                dvt0w = 0                         
+       dvt1w = 0                                dvt2w = 0                                 dsub = 0.1                               minv = 0.05                      
+       voffl = 0                                dvtp0 = 1.000e-10                        dvtp1 = 0.1                               lpe0 = 0                         
+        lpeb = 0                                ngate = 3.000e+20                          nsd = 2.000e+20                         phin = 0                         
+        cdsc = 0                                cdscb = 0                                cdscd = 0                                  cit = 0                         
+        voff = {AGAUSS(-0.13, 0.00650, 1)}        etab = 0                                  vfb = -0.55                               ua = 6.000e-10                 
+          ub = 1.200e-18                           uc = 0                                   a0 = 1                                  ags = 0                         
+          a1 = 0                                   a2 = 1                                   b0 = 0                                   b1 = 0                         
+        keta = 0.04                               dwg = 0                                  dwb = 0                                 pclm = 0.02                      
+     pdiblc1 = 0.001                          pdiblc2 = 0.001                          pdiblcb = -0.005                           drout = 0.5                       
+        pvag = 1.000e-20                        delta = 0.01                            pscbe1 = 8.140e+08                       pscbe2 = 1.000e-07                 
+      fprout = 0.2                              pdits = 0.08                            pditsd = 0.23                            pditsl = 2300000                   
+         rsh = 5                                  rsw = 80                                 rdw = 80                             rdswmin = 0                         
+      rdwmin = 0                               rswmin = 0                                 prwg = 0                                 prwb = 0                         
+          wr = 1                               alpha0 = 0.074                           alpha1 = 0.005                            beta0 = 30                        
+       agidl = 2.000e-04                        bgidl = 2.100e+09                        cgidl = 2.000e-04                        egidl = 0.8                       
+     aigbacc = 0.012                          bigbacc = 0.0028                         cigbacc = 0.002                          nigbacc = 1                         
+     aigbinv = 0.014                          bigbinv = 0.004                          cigbinv = 0.004                          eigbinv = 1.1                       
+     nigbinv = 3                                 aigc = 0.02                              bigc = 0.0027                            cigc = 0.002                     
+       aigsd = 0.02                             bigsd = 0.0027                           cigsd = 0.002                             nigc = 1                         
+     poxedge = 1                                pigcd = 1                                 ntox = 1                               xrcrg1 = 12                        
+      xrcrg2 = 5                                 cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                 
+     ckappas = 0.03                           ckappad = 0.03                              acde = 1                                 moin = 15                        
+        noff = 0.9                             voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                         
+         kt2 = 0.022                              ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                 
+         uc1 = -5.600e-11                         prt = 0                                   at = 33000                          fnoimod = 1                         
+     tnoimod = 0                                  jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                 
+         njs = 1                             ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                        
+       xjbvs = 1                                  jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                 
+         njd = 1                             ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                        
+       xjbvd = 1                                  pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                       
+       pbsws = 1                                cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                         
+      cjswgs = 3.000e-10                       mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                 
+         mjd = 0.5                              pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                      
+      pbswgd = 1                               cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                     
+         tcj = 0.001                            tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                     
+      tcjswg = 0.001                             xtis = 3                                 xtid = 3                                 dmcg = 0                         
+        dmci = 0                                 dmdg = 0                                dmcgt = 0                                  dwj = 0                         
+         xgw = 0                                  xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                 
+        rbpb = 5                                 rbpd = 15                                rbps = 15                                rbdb = 15                        
+        rbsb = 15                               ngcon = 1                         

.model  NMOS_VTH  nmos
+       level = 54                                tnom = 27                              epsrox = 3.9                               eta0 = 0.008                     
+     nfactor = 1.6                               wint = 5.000e-09                         cgso = 1.100e-10                         cgdo = 1.100e-10                 
+        toxe = 1.630e-09                         toxp = 1.000e-09                         toxm = 1.630e-09                       toxref = 1.630e-09                 
+        dtox = 6.300e-10                         lint = 3.750e-09                         vth0 = {AGAUSS(0.6078, 0.03039, 1)}          k1 = 0.4                       
+          u0 = {AGAUSS(0.049, 0.00245, 1)}        vsat = 170000                            rdsw = 155                               ndep = 3.240e+18                 
+          xj = 1.980e-08                      version = 4.8                            binunit = 1                             paramchk = 1                         
+      mobmod = 0                               capmod = 2                               igcmod = 1                               igbmod = 1                         
+      geomod = 1                               diomod = 1                               rdsmod = 0                             rbodymod = 1                         
+    rgatemod = 1                               permod = 1                             acnqsmod = 0                             trnqsmod = 0                         
+          ll = 0                                   wl = 0                                  lln = 1                                  wln = 1                         
+          lw = 0                                   ww = 0                                  lwn = 1                                  wwn = 1                         
+         lwl = 0                                  wwl = 0                                xpart = 0                                   k2 = 0                         
+          k3 = 0                                  k3b = 0                                   w0 = 2.500e-06                         dvt0 = 1                         
+        dvt1 = 2                                 dvt2 = 0                                dvt0w = 0                                dvt1w = 0                         
+       dvt2w = 0                                 dsub = 0.1                               minv = 0.05                             voffl = 0                         
+       dvtp0 = 1.000e-10                        dvtp1 = 0.1                               lpe0 = 0                                 lpeb = 0                         
+       ngate = 3.000e+20                          nsd = 2.000e+20                         phin = 0                                 cdsc = 0                         
+       cdscb = 0                                cdscd = 0                                  cit = 0                                 voff = {AGAUSS(-0.13, 0.00650, 1)}
+        etab = 0                                  vfb = -0.55                               ua = 6.000e-10                           ub = 1.200e-18                 
+          uc = 0                                   a0 = 1                                  ags = 0                                   a1 = 0                         
+          a2 = 1                                   b0 = 0                                   b1 = 0                                 keta = 0.04                      
+         dwg = 0                                  dwb = 0                                 pclm = 0.02                           pdiblc1 = 0.001                     
+     pdiblc2 = 0.001                          pdiblcb = -0.005                           drout = 0.5                               pvag = 1.000e-20                 
+       delta = 0.01                            pscbe1 = 8.140e+08                       pscbe2 = 1.000e-07                       fprout = 0.2                       
+       pdits = 0.08                            pditsd = 0.23                            pditsl = 2300000                            rsh = 5                         
+         rsw = 80                                 rdw = 80                             rdswmin = 0                               rdwmin = 0                         
+      rswmin = 0                                 prwg = 0                                 prwb = 0                                   wr = 1                         
+      alpha0 = 0.074                           alpha1 = 0.005                            beta0 = 30                               agidl = 2.000e-04                 
+       bgidl = 2.100e+09                        cgidl = 2.000e-04                        egidl = 0.8                            aigbacc = 0.012                     
+     bigbacc = 0.0028                         cigbacc = 0.002                          nigbacc = 1                              aigbinv = 0.014                     
+     bigbinv = 0.004                          cigbinv = 0.004                          eigbinv = 1.1                            nigbinv = 3                         
+        aigc = 0.015211                          bigc = 0.0027432                         cigc = 0.002                            aigsd = 0.015211                  
+       bigsd = 0.0027432                        cigsd = 0.002                             nigc = 1                              poxedge = 1                         
+       pigcd = 1                                 ntox = 1                               xrcrg1 = 12                              xrcrg2 = 5                         
+        cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                      ckappas = 0.03                      
+     ckappad = 0.03                              acde = 1                                 moin = 15                                noff = 0.9                       
+      voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                                  kt2 = 0.022                     
+         ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                          uc1 = -5.600e-11                
+         prt = 0                                   at = 33000                          fnoimod = 1                              tnoimod = 0                         
+         jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                          njs = 1                         
+    ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                               xjbvs = 1                         
+         jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                          njd = 1                         
+    ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                               xjbvd = 1                         
+         pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                              pbsws = 1                         
+       cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                               cjswgs = 3.000e-10                 
+      mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                          mjd = 0.5                       
+       pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                            pbswgd = 1                         
+      cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                              tcj = 0.001                     
+       tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                           tcjswg = 0.001                     
+        xtis = 3                                 xtid = 3                                 dmcg = 0                                 dmci = 0                         
+        dmdg = 0                                dmcgt = 0                                  dwj = 0                                  xgw = 0                         
+         xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                         rbpb = 5                         
+        rbpd = 15                                rbps = 15                                rbdb = 15                                rbsb = 15                        
+       ngcon = 1                         

.model  PMOS_VTH  pmos
+       level = 54                             version = 4.8                            binunit = 1                             paramchk = 1                         
+      mobmod = 0                               capmod = 2                               igcmod = 1                               igbmod = 1                         
+      geomod = 1                               diomod = 1                               rdsmod = 0                             rbodymod = 1                         
+    rgatemod = 1                               permod = 1                             acnqsmod = 0                             trnqsmod = 0                         
+        tnom = 27                                toxe = 1.600e-09                         toxp = 1.000e-09                         toxm = 1.600e-09                 
+        dtox = 6.000e-10                       epsrox = 3.9                               wint = 5.000e-09                         lint = 3.750e-09                 
+          ll = 0                                   wl = 0                                  lln = 1                                  wln = 1                         
+          lw = 0                                   ww = 0                                  lwn = 1                                  wwn = 1                         
+         lwl = 0                                  wwl = 0                                xpart = 0                               toxref = 1.600e-09                 
+        vth0 = {AGAUSS(-0.5044, 0.02522, 1)}          k1 = 0.4                                 k2 = -0.01                               k3 = 0                         
+         k3b = 0                                   w0 = 2.500e-06                         dvt0 = 1                                 dvt1 = 2                         
+        dvt2 = -0.032                           dvt0w = 0                                dvt1w = 0                                dvt2w = 0                         
+        dsub = 0.1                               minv = 0.05                             voffl = 0                                dvtp0 = 1.000e-11                 
+       dvtp1 = 0.05                              lpe0 = 0                                 lpeb = 0                                   xj = 1.400e-08                 
+       ngate = 2.000e+20                         ndep = 2.440e+18                          nsd = 2.000e+20                         phin = 0                         
+        cdsc = 0                                cdscb = 0                                cdscd = 0                                  cit = 0                         
+        voff = {AGAUSS(-0.126, 0.00630, 1)}     nfactor = 1.8                               eta0 = 0.0125                            etab = 0                         
+         vfb = 0.55                                u0 = {AGAUSS(0.021, 0.00105, 1)}          ua = 2.000e-09                           ub = 5.000e-19                 
+          uc = 0                                 vsat = 80000                               a0 = 1                                  ags = 1.000e-20                 
+          a1 = 0                                   a2 = 1                                   b0 = 0                                   b1 = 0                         
+        keta = -0.047                             dwg = 0                                  dwb = 0                                 pclm = 0.12                      
+     pdiblc1 = 0.001                          pdiblc2 = 0.001                          pdiblcb = 3.400e-08                        drout = 0.56                      
+        pvag = 1.000e-20                        delta = 0.01                            pscbe1 = 8.140e+08                       pscbe2 = 9.580e-07                 
+      fprout = 0.2                              pdits = 0.08                            pditsd = 0.23                            pditsl = 2300000                   
+         rsh = 5                                 rdsw = 250                                rsw = 75                                 rdw = 75                        
+     rdswmin = 0                               rdwmin = 0                               rswmin = 0                                 prwg = 0                         
+        prwb = 0                                   wr = 1                               alpha0 = 0.074                           alpha1 = 0.005                     
+       beta0 = 30                               agidl = 2.000e-04                        bgidl = 2.100e+09                        cgidl = 2.000e-04                 
+       egidl = 0.8                            aigbacc = 0.012                          bigbacc = 0.0028                         cigbacc = 0.002                     
+     nigbacc = 1                              aigbinv = 0.014                          bigbinv = 0.004                          cigbinv = 0.004                     
+     eigbinv = 1.1                            nigbinv = 3                                 aigc = 0.0097                            bigc = 0.00125                   
+        cigc = 8.000e-04                        aigsd = 0.0097                           bigsd = 0.00125                          cigsd = 8.000e-04                 
+        nigc = 1                              poxedge = 1                                pigcd = 1                                 ntox = 1                         
+      xrcrg1 = 12                              xrcrg2 = 5                                 cgso = 1.100e-10                         cgdo = 1.100e-10                 
+        cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                      ckappas = 0.03                      
+     ckappad = 0.03                              acde = 1                                 moin = 15                                noff = 0.9                       
+      voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                                  kt2 = 0.022                     
+         ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                          uc1 = -5.600e-11                
+         prt = 0                                   at = 33000                          fnoimod = 1                              tnoimod = 0                         
+         jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                          njs = 1                         
+    ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                               xjbvs = 1                         
+         jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                          njd = 1                         
+    ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                               xjbvd = 1                         
+         pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                              pbsws = 1                         
+       cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                               cjswgs = 3.000e-10                 
+      mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                          mjd = 0.5                       
+       pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                            pbswgd = 1                         
+      cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                              tcj = 0.001                     
+       tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                           tcjswg = 0.001                     
+        xtis = 3                                 xtid = 3                                 dmcg = 0                                 dmci = 0                         
+        dmdg = 0                                dmcgt = 0                                  dwj = 0                                  xgw = 0                         
+         xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                         rbpb = 5                         
+        rbpd = 15                                rbps = 15                                rbdb = 15                                rbsb = 15                        
+       ngcon = 1                         

.model  PMOS_VTG  pmos
+       level = 54                                vth0 = {AGAUSS(-0.3842, 0.01921, 1)}      toxref = 1.260e-09                         vsat = 62000                     
+        toxe = 1.260e-09                         toxp = 1.000e-09                         toxm = 1.260e-09                         dtox = 2.600e-10                 
+      epsrox = 3.9                               wint = 5.000e-09                         lint = 3.750e-09                      version = 4.8                       
+     binunit = 1                             paramchk = 1                               mobmod = 0                               capmod = 2                         
+      igcmod = 1                               igbmod = 1                               geomod = 1                               diomod = 1                         
+      rdsmod = 0                             rbodymod = 1                             rgatemod = 1                               permod = 1                         
+    acnqsmod = 0                             trnqsmod = 0                                 tnom = 27                                  ll = 0                         
+          wl = 0                                  lln = 1                                  wln = 1                                   lw = 0                         
+          ww = 0                                  lwn = 1                                  wwn = 1                                  lwl = 0                         
+         wwl = 0                                xpart = 0                                   xl = -2.000e-08                          k1 = 0.4                       
+          k2 = -0.01                               k3 = 0                                  k3b = 0                                   w0 = 2.500e-06                 
+        dvt0 = 1                                 dvt1 = 2                                 dvt2 = -0.032                           dvt0w = 0                         
+       dvt1w = 0                                dvt2w = 0                                 dsub = 0.1                               minv = 0.05                      
+       voffl = 0                                dvtp0 = 1.000e-11                        dvtp1 = 0.05                              lpe0 = 0                         
+        lpeb = 0                                   xj = 1.980e-08                        ngate = 2.000e+20                         ndep = 2.440e+18                 
+         nsd = 2.000e+20                         phin = 0                                 cdsc = 0                                cdscb = 0                         
+       cdscd = 0                                  cit = 0                                 voff = {AGAUSS(-0.126, 0.00630, 1)}     nfactor = 2.22                      
+        eta0 = 0.0055                            etab = 0                                  vfb = 0.55                                u0 = {AGAUSS(0.02, 0.00100, 1)}
+          ua = 2.000e-09                           ub = 5.000e-19                           uc = 0                                   a0 = 1                         
+         ags = 1.000e-20                           a1 = 0                                   a2 = 1                                   b0 = 0                         
+          b1 = 0                                 keta = -0.047                             dwg = 0                                  dwb = 0                         
+        pclm = 0.12                           pdiblc1 = 0.001                          pdiblc2 = 0.001                          pdiblcb = 3.400e-08                 
+       drout = 0.56                              pvag = 1.000e-20                        delta = 0.01                            pscbe1 = 8.140e+08                 
+      pscbe2 = 9.580e-07                       fprout = 0.2                              pdits = 0.08                            pditsd = 0.23                      
+      pditsl = 2300000                            rsh = 5                                 rdsw = 155                                rsw = 75                        
+         rdw = 75                             rdswmin = 0                               rdwmin = 0                               rswmin = 0                         
+        prwg = 0                                 prwb = 0                                   wr = 1                               alpha0 = 0.074                     
+      alpha1 = 0.005                            beta0 = 30                               agidl = 2.000e-04                        bgidl = 2.100e+09                 
+       cgidl = 2.000e-04                        egidl = 0.8                            aigbacc = 0.012                          bigbacc = 0.0028                    
+     cigbacc = 0.002                          nigbacc = 1                              aigbinv = 0.014                          bigbinv = 0.004                     
+     cigbinv = 0.004                          eigbinv = 1.1                            nigbinv = 3                                 aigc = 0.010687                  
+        bigc = 0.0012607                         cigc = 8.000e-04                        aigsd = 0.010687                         bigsd = 0.0012607                 
+       cigsd = 8.000e-04                         nigc = 1                              poxedge = 1                                pigcd = 1                         
+        ntox = 1                               xrcrg1 = 12                              xrcrg2 = 5                                 cgso = 1.100e-10                 
+        cgdo = 1.100e-10                         cgbo = 2.560e-11                         cgdl = 2.653e-10                         cgsl = 2.653e-10                 
+     ckappas = 0.03                           ckappad = 0.03                              acde = 1                                 moin = 15                        
+        noff = 0.9                             voffcv = 0.02                               kt1 = -0.11                             kt1l = 0                         
+         kt2 = 0.022                              ute = -1.5                               ua1 = 4.310e-09                          ub1 = 7.610e-18                 
+         uc1 = -5.600e-11                         prt = 0                                   at = 33000                          fnoimod = 1                         
+     tnoimod = 0                                  jss = 1.000e-04                         jsws = 1.000e-11                        jswgs = 1.000e-10                 
+         njs = 1                             ijthsfwd = 0.01                          ijthsrev = 0.001                              bvs = 10                        
+       xjbvs = 1                                  jsd = 1.000e-04                         jswd = 1.000e-11                        jswgd = 1.000e-10                 
+         njd = 1                             ijthdfwd = 0.01                          ijthdrev = 0.001                              bvd = 10                        
+       xjbvd = 1                                  pbs = 1                                  cjs = 5.000e-04                          mjs = 0.5                       
+       pbsws = 1                                cjsws = 5.000e-10                        mjsws = 0.33                            pbswgs = 1                         
+      cjswgs = 3.000e-10                       mjswgs = 0.33                               pbd = 1                                  cjd = 5.000e-04                 
+         mjd = 0.5                              pbswd = 1                                cjswd = 5.000e-10                        mjswd = 0.33                      
+      pbswgd = 1                               cjswgd = 5.000e-10                       mjswgd = 0.33                               tpb = 0.005                     
+         tcj = 0.001                            tpbsw = 0.005                            tcjsw = 0.001                           tpbswg = 0.005                     
+      tcjswg = 0.001                             xtis = 3                                 xtid = 3                                 dmcg = 0                         
+        dmci = 0                                 dmdg = 0                                dmcgt = 0                                  dwj = 0                         
+         xgw = 0                                  xgl = 0                                 rshg = 0.4                              gbmin = 1.000e-10                 
+        rbpb = 5                                 rbpd = 15                                rbps = 15                                rbdb = 15                        
+        rbsb = 15                        


